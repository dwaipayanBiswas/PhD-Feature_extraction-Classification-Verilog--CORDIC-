//*********************************************************************************************
// Test Bench
// Author: Dwaipayan Biswas
// Email: db9g10@ecs.soton.ac.uk
// University of Southampton
//*********************************************************************************************
`timescale 1ns / 100ps
`include "parameter.v"

module feature_select_stim;

parameter period = 100000;

reg [15:0] dataIn;
reg clk, nReset, nRd, nWr, nCs;
reg [2:0] Addr;

wire [15:0] dataOut;
wire Intr; 

feature_select dut (clk, nReset, Addr, dataIn, dataOut, nRd, nWr, nCs, Intr);

task wr_data;
input [2:0] address;
input [15:0] data;
	begin
	#period
	Addr = address;
	dataIn = data;
	nCs = 0;
	nRd = 1;
	nWr = 0;
#period;
Addr = address;
dataIn = 16'bZ;
nCs = 1;
nRd = 1;
nWr = 1;
#period;
end
endtask

task rd_data;
input [2:0] address;
begin
#period;
Addr = address;
nCs = 0;
nRd = 0;
nWr = 1;
#period;
Addr = address;
nCs = 1;
nRd = 1;
nWr = 1;
#period;
end
endtask

always
begin
  clk = 1;
  #(period/2)	clk = 0;
  #(period/2)	clk = 1;
end


initial
begin
nReset= 0; 
dataIn = 16'bZ;
Addr = 3'b000;
nRd = 1;
nWr = 1;
nCs = 1;		 
#(10*period);
nReset= 1;
#(20*period);
// write feature code
wr_data (3'b110,16'b0000011011110000);
wr_data (3'b111, 16'b0000000011111110);
rd_data (3'b110);
rd_data (3'b111);	    
// write start, select X
wr_data (3'b010,16'h8000);
rd_data (3'b010);
#(20*period);

// x data
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);

#(2000*period);

// remove start, select y, write start
wr_data (3'b010,16'h0001);
#(20*period);
wr_data (3'b010,16'h8001);
#(20*period);



// y data
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000010000);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001110);
#(2*period); wr_data(3'b000,16'b0000000000001111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);

#(2000*period);

// remove start, select z, write start
wr_data (3'b010,16'h0003);
#(20*period);
wr_data (3'b010,16'h8003);
#(20*period);

// z data

#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001100);
#(2*period); wr_data(3'b000,16'b0000000000001101);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001011);
#(2*period); wr_data(3'b000,16'b0000000000001001);
#(2*period); wr_data(3'b000,16'b0000000000001010);
#(2*period); wr_data(3'b000,16'b0000000000001000);
#(2*period); wr_data(3'b000,16'b0000000000000111);
#(2*period); wr_data(3'b000,16'b0000000000001101);

#(2000*period);

// remove start, select z, write start
wr_data (3'b010,16'h0000);
#(20*period);
wr_data (3'b010,16'h8000);
#(20*period);

// x cent
#(2*period); wr_data(3'b001,16'b0000000000001011);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001010);
#(2*period); wr_data(3'b001,16'b0000000000001011);
#(2*period); wr_data(3'b001,16'b0000000000001010);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001010);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001010);

// y cent

#(2000*period);

// remove start, select z, write start
wr_data (3'b010,16'h0001);
#(20*period);
wr_data (3'b010,16'h8001);
#(20*period);

#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000010000);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001110);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000010000);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001111);
#(2*period); wr_data(3'b001,16'b0000000000001110);

// z cent

#(2000*period);

// remove start, select z, write start
wr_data (3'b010,16'h0007);
#(20*period);
wr_data (3'b010,16'h8007);
#(20*period);

#(2*period); wr_data(3'b001,16'b0000000000001010);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001001);
#(2*period); wr_data(3'b001,16'b0000000000001000);
#(2*period); wr_data(3'b001,16'b0000000000001011);
#(2*period); wr_data(3'b001,16'b0000000000001011);
#(2*period); wr_data(3'b001,16'b0000000000001001);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001000);
#(2*period); wr_data(3'b001,16'b0000000000001000);
#(2*period); wr_data(3'b001,16'b0000000000000111);
#(2*period); wr_data(3'b001,16'b0000000000001011);
#(2*period); wr_data(3'b001,16'b0000000000001000);
#(2*period); wr_data(3'b001,16'b0000000000001001);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000001010);
#(2*period); wr_data(3'b001,16'b0000000000001001);
#(2*period); wr_data(3'b001,16'b0000000000001000);
#(2*period); wr_data(3'b001,16'b0000000000001010);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001000);
#(2*period); wr_data(3'b001,16'b0000000000001010);
#(2*period); wr_data(3'b001,16'b0000000000001100);
#(2*period); wr_data(3'b001,16'b0000000000000111);
#(2*period); wr_data(3'b001,16'b0000000000001011);
#(2*period); wr_data(3'b001,16'b0000000000001101);
#(2*period); wr_data(3'b001,16'b0000000000001001);
#(2*period); wr_data(3'b001,16'b0000000000001000);


#(1000*period);

rd_data (3'b000);
rd_data (3'b001);
rd_data (3'b010);
rd_data (3'b011);
rd_data (3'b100);
rd_data (3'b101);
rd_data (3'b110);
rd_data (3'b111);

#(10*period);

end

endmodule
